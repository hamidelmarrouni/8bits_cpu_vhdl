library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;
use std.textio.all;
use work.constants_pkg.all;

entity memory is
  generic (
    MEM_SIZE  : natural := MEM_SIZE_C;     -- e.g. 4096 bytes
    INIT_FILE : string  := "program.hex"   -- used ONLY IN SIMULATION
  );
  port (
    clk   : in  std_logic;
    addr  : in  std_logic_vector(ADDR_W-1 downto 0);
    dout  : in  std_logic_vector(DATA_W-1 downto 0); -- data from CPU to write
    din   : out std_logic_vector(DATA_W-1 downto 0); -- data to CPU
    rd    : in  std_logic;
    wr    : in  std_logic;
    ready : out std_logic
  );
end entity;

architecture rtl of memory is

  ----------------------------------------------------------------------
  -- MEMORY ARRAY DECLARATION
  ----------------------------------------------------------------------
  type mem_t is array (0 to MEM_SIZE-1) of std_logic_vector(DATA_W-1 downto 0);

  ----------------------------------------------------------------------
  -- SIMULATION-ONLY INITIALIZATION (READ program.hex)
  --
  -- This part uses file I/O ? NOT SYNTHESIZABLE.
  -- It is wrapped inside synthesis translate_off/on so FPGA tools ignore it.
  --
  -- REAL HARDWARE:
  --   Memory starts empty and is filled by the UART bootloader.
  --
  -- SIMULATION:
  --   Memory is initialized from program.hex generated by Python GUI.
  ----------------------------------------------------------------------
  -- synthesis translate_off
  impure function init_mem(fname : in string) return mem_t is
    file     f      : text open read_mode is fname;
    variable l      : line;
    variable m      : mem_t := (others => (others => '0'));
    variable idx    : integer := 0;
    variable data_v : std_logic_vector(DATA_W-1 downto 0);
  begin
    if fname'length = 0 then
      return m;  -- no init file ? memory all zeros
    end if;

    -- Read 1 byte per line (2 hex characters)
    while not endfile(f) and idx < MEM_SIZE loop
      readline(f, l);
      if l'length > 0 then
        hread(l, data_v);
        m(idx) := data_v;
        idx    := idx + 1;
      end if;
    end loop;

    return m;
  end function;
  -- synthesis translate_on

  ----------------------------------------------------------------------
  -- MEMORY SIGNAL
  --
  -- SIMULATION:
  --     initialized using init_mem(INIT_FILE)
  --
  -- REAL FPGA:
  --     synthesis will IGNORE init_mem ? memory starts empty (all zeros)
  --     UART loader will write program into memory at runtime
  ----------------------------------------------------------------------
  signal mem : mem_t :=
  -- synthesis translate_off
      init_mem(INIT_FILE)
  -- synthesis translate_on
  -- synthesis translate_off
  ;
  -- synthesis translate_on

  signal rdata_reg : std_logic_vector(DATA_W-1 downto 0) := (others => '0');

  -- address integer
  signal addr_i : integer range 0 to MEM_SIZE-1;

begin

  ----------------------------------------------------------------------
  -- ADDRESS DECODE
  ----------------------------------------------------------------------
  addr_i <= to_integer(unsigned(addr));

  ----------------------------------------------------------------------
  -- SYNCHRONOUS READ/WRITE (1-cycle read latency)
  ----------------------------------------------------------------------
  process(clk)
  begin
    if rising_edge(clk) then

      ------------------------------------------------------------------
      -- WRITE OPERATION
      --
      -- In REAL FPGA: written by CPU or UART bootloader
      -- In SIMULATION: same behavior
      ------------------------------------------------------------------
      if wr = '1' then
        if addr_i < MEM_SIZE then
          mem(addr_i) <= dout;
        end if;
      end if;

      ------------------------------------------------------------------
      -- READ OPERATION (REGISTERED, 1-cycle latency)
      ------------------------------------------------------------------
      if rd = '1' then
        if addr_i < MEM_SIZE then
          rdata_reg <= mem(addr_i);
        else
          rdata_reg <= (others => '0');
        end if;
      end if;

    end if;
  end process;

  din   <= rdata_reg;

  ----------------------------------------------------------------------
  -- ALWAYS READY (no wait states)
  -- Compatible with your simple CPU design
  ----------------------------------------------------------------------
  ready <= '1';

end architecture;
